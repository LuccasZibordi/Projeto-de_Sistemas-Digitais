LIBRARY ieee;
use ieee.std_logic_1164.all;
use work.all;

entity comparador is
port( x,y: in std_logic_vector (3 downto 0);
AeqB, AgtB,AltB: out std_logic);
end comparador;

Architecture compare of comparador is
signal i: std_logic_vector (3 downto 0);
signal eq,gr: std_logic;

begin
i(3) <= x(0) xnor y(0);
i(2) <= x(1) xnor y(1);
i(1) <= x(2) xnor y(2);
i(0) <= x(3) xnor y(3);

eq <= i(0) and i(1) and  i(2) and i(3);
gr <= (x(3) and not y(3)) or (i(3) and x(2) and not y(2)) or (i(2) and i(3) and x(1) and not y(1)) or (i(1) and i(2) and i(3) and x(0) and not y(0));
AeqB <= eq;
AgtB <= gr;
AltB <= eq nor gr;
end compare;